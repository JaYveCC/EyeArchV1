`define PORT_EXPONENT 3 //amount of ports = 2^PORT_EXPONENT
