`define PORT_EXPONENT 1 //amount of ports = 2^PORT_EXPONENT
