`define PORT_EXPONENT 3 //anmount of ports = 2^PORT_EXPONENT
